module hitsz
endmodule
