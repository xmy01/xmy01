module hitsz
  sbxiantao
endmodule
