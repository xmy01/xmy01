module hitwh
endmodule
