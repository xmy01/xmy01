module hitwh
  hitwh
endmodule
