module hitsz
  sbhitwh
endmodule
